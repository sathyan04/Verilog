module sub(input [3:0]a,b, output [4:0]diff);
assign diff=a-b;
endmodule
