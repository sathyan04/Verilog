module sr_latch(input s,r, output reg q);
always @(*) begin
	if(s==1'b0 && r==1'b1)
		q=1'b0;
	else if (s==1'b1 && r==1'b0) 
		q=1'b1;
	else if (s==1'b1 && r==1'b1)
		q=1'bx;
end
endmodule
