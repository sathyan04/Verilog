`default_nettype none
module top_module(
    input a,
    input b,
    input c,
    input d,
    output out,
    output out_n   ); 
	wire x,y,z;
    and(x,a,b);
    and(y,c,d);
    or(z,x,y);
    assign out=z;
    not(out_n,out);
endmodule
