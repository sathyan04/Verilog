module mul(input [3:0]a,b, output [7:0]m);
assign m=a*b;
endmodule
