module natural(input [3:0]n, output [3:0]sum);
assign sum=(n*(n+1))/2;
endmodule

