module btxs(input [3:0]bin, output [3:0]exs);
assign exs = bin + 4'b0011;
endmodule

