module sequence_detector_1101_tb();
reg clk,rst,data;
reg [1:0] mode;
wire detected;
sequence_detector_1101 dut(.clk(clk),.rst(rst),.data(data),.mode(mode),.detected(detected));
initial begin
	clk=0;
	forever #5 clk=~clk;
end
initial begin
	$dumpfile("sequencegtk.vcd");
	$dumpvars(0);
	rst=1;data=0;#10;rst=0;
	$display("Moore Overlap");
	mode=2'b00;
	data=1;#10;
	data=1;#10;
	data=0;#10;
	data=1;#10;
	data=1;#10;
        data=0;#10;
	data=1;#10;
	data=1;#10;
        data=0;#10;
	data=1;#10;
	data=1;#10;
        data=0;#10;
	data=1;#10;
	data=1;#10;
        data=0;#10;
	data=1;#10;
	data=1;#10;
        data=0;#30;
	$display("\nMoore Non Overlap");
	mode=2'b01;
	data=1;#10;
        data=1;#10;
        data=0;#10;
	data=1;#10;
        data=1;#10;
        data=0;#10;
	data=1;#10;
        data=1;#10;
        data=0;#10;
	data=1;#10;
        data=1;#10;
        data=0;#10;
	data=1;#10;
        data=1;#10;
        data=0;#10;
	data=1;#10;
        data=1;#10;
        data=0;#30;
	$display("\nMealy Overlap");
	mode=2'b10;
        data=1;#10;
	data=1;#10;
        data=0;#10;
        data=1;#10;
	data=1;#10;
        data=0;#10;
        data=1;#10;
	data=1;#10;
        data=0;#10;
        data=1;#10;
	data=1;#10;
        data=0;#10;
        data=1;#10;
	data=1;#10;
        data=0;#10;
        data=1;#10;
	data=1;#10;
        data=0;#30;
	$display("\nMealy Non Overlap");
	mode=2'b11;
	data=1;#10;
        data=1;#10;
        data=0;#10;
	data=1;#10;
        data=1;#10;
        data=0;#10;
	data=1;#10;
        data=1;#10;
        data=0;#10;
	data=1;#10;
        data=1;#10;
        data=0;#10;
	data=1;#10;
        data=1;#10;
        data=0;#10;
	data=1;#10;
        data=1;#10;
        data=0;#10;
	$finish;
end
always@(posedge clk) begin
	if(!rst)
		$display("Data=%b | Output=%b",data, detected);
end
endmodule
